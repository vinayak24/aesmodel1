module Inv_Round_Last(Clk,RIn,KeyIn,Out);
  input Clk;
  input [127:0]RIn;
  input [127:0]KeyIn;
  output [127:0]Out;
  wire [127:0] ISubBytes,ISR;
  
//  KeyGeneration M0(Round_Count,KeyLastIn,Key_Out);


  Inv_ShiftRow M2(RIn,ISR);
  Inv_SubBytes M1(ISR,ISubBytes);  
  assign Out= KeyIn^ISubBytes;
  
endmodule