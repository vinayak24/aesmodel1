module Inv_ShiftRow (In,Out);
  input [127:0]In;
  output [127:0]Out;
  assign Out[127:120] = In[127:120];
  assign Out[119:112] = In[23:16];
  assign Out[111:104] = In[47:40];
  assign Out[103:96]  = In[71:64];
  assign Out[95:88]   = In[95:88];
  assign Out[87:80]   = In[119:112];
  assign Out[79:72]   = In[15:8];
  assign Out[71:64]   = In[39:32];
  assign Out[63:56]   = In[63:56];
  assign Out[55:48]   = In[87:80];
  assign Out[47:40]   = In[111:104];
  assign Out[39:32]   = In[7:0];
  assign Out[31:24]   = In[31:24];
  assign Out[23:16]   = In[55:48];
  assign Out[15:8]    = In[79:72];
  assign Out[7:0]     = In[103:96];
  
endmodule